Library ieee;
use ieee.std_logic_1164.all;

ENTITY unidade_contole IS
	PORT(OPCode: IN STD_LOGIC_VECTOR (5 DOWNTO 0);
		  